module adder (
    input a, 
    input b,
    output sum,
);
    assign sum = a+b;
    
endmodule